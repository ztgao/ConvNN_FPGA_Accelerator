// version 1.0 -- setup
// Description:
// For a better view of IEEE-754 format.

module type_cast(



);

// $bitstoshortreal