// version 1.0 -- 	12.09
//					setup
// Description:

`include "../../global_define.v"
module conv_layer_output_interface(	
//--input
	clk,
	rst_n,
	data_in,
	valid_in,
//--output
	data_out
);

